package Accelerator;
	import Defines::*;

	interface Ifc_Accelerator;
		interface MemClient portA;
		interface MemClient portB;
	endinterface

endpackage
